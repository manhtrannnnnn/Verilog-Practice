//---------------------------------------- 8x8 sequential multiplexer ----------------------------------------//

module seq_multiplexer(
    input clk,
    input asyn_reset,
    input syn_load,
    input [7:0] a,
    input [7:0] b,
    output [15:0] result,
    output valid
);
endmodule