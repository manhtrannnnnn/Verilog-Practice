//-----------------------------------------------Design 16 x 16 bidirectional memory-----------------------------------------------//
module bidirectional_mem();

endmodule