//----------------------------------- Parity Generator -----------------------------------//
module parity(
    input clk, asyn_rst,
    input valid_in,
    input data_in,
    output 
):
endmodule