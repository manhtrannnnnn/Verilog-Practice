//---------------------------------------- 8x8 sequential multiplexer ----------------------------------------//

module seq_multiplexer(
    input rst_n, syn_load, 
    output valid
);
endmodule